module clk(clock);

input clock;

endmodule